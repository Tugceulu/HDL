//////////////////////////////////////////////////////////////////////////////
//Alwaysblock1(combinational)
//Combinational: always @(*)
//Clocked: always @(posedge clk)
//assign out1 = a & b | c ^ d;
//always @(*) out2 = a & b | c ^ d;
// synthesis verilog_input_version verilog_2001
module top_module(
    input a, 
    input b,
    output wire out_assign,
    output reg out_alwaysblock
);
 	assign out_assign = a & b;
    always @(*) begin
        out_alwaysblock = a & b;
    end
endmodule

//////////////////////////////////////////////////////////////////////////////
//Alwaysblock2(closed)

//////////////////////////////////////////////////////////////////////////////
//If statement

//////////////////////////////////////////////////////////////////////////////
//If statement latches

//////////////////////////////////////////////////////////////////////////////
//Case statement

//////////////////////////////////////////////////////////////////////////////
//Priority encoder

//////////////////////////////////////////////////////////////////////////////
//Priority encoder with casez

//////////////////////////////////////////////////////////////////////////////
//Avoiding latches

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//
