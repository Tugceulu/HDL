//////////////////////////////////////////////////////////////////////////////
//Alwaysblock1(combinational)
//Combinational: always @(*)
//Clocked: always @(posedge clk)
//assign out1 = a & b | c ^ d;
//always @(*) out2 = a & b | c ^ d;
// synthesis verilog_input_version verilog_2001
module top_module(
    input a, 
    input b,
    output wire out_assign,
    output reg out_alwaysblock
);
 	assign out_assign = a & b;
    always @(*) begin
        out_alwaysblock = a & b;
    end
endmodule

//////////////////////////////////////////////////////////////////////////////
//Alwaysblock2(closed)
// synthesis verilog_input_version verilog_2001
module top_module(
    input clk,
    input a,
    input b,
    output wire out_assign,
    output reg out_always_comb,
    output reg out_always_ff   );
    
	assign out_assign=a^b;
    always @(*) begin
        out_always_comb=a^b;
    end
    always @(posedge clk) begin
        out_always_ff=a^b;
    end
endmodule

//////////////////////////////////////////////////////////////////////////////
//If statement
// synthesis verilog_input_version verilog_2001
module top_module(
    input a,
    input b,
    input sel_b1,
    input sel_b2,
    output wire out_assign,
    output reg out_always   ); 
	
    always @(*) begin
        case(sel_b1&sel_b2)
            0:out_always=a;
            1:out_always=b;
        endcase
    end        
    assign out_assign= out_always;
endmodule

//////////////////////////////////////////////////////////////////////////////
//If statement latches
// synthesis verilog_input_version verilog_2001
module top_module (
    input      cpu_overheated,
    output reg shut_off_computer,
    input      arrived,
    input      gas_tank_empty,
    output reg keep_driving  ); //
	always @(*) begin
        if (cpu_overheated)
           shut_off_computer = 1;
        else
            shut_off_computer = 0;
    end

    always @(*) begin
        if (~arrived)
           keep_driving = ~gas_tank_empty;
        else 
            keep_driving=0;          
    end
endmodule

//////////////////////////////////////////////////////////////////////////////
//Case statement
// synthesis verilog_input_version verilog_2001
module top_module ( 
    input [2:0] sel, 
    input [3:0] data0,
    input [3:0] data1,
    input [3:0] data2,
    input [3:0] data3,
    input [3:0] data4,
    input [3:0] data5,
    output reg [3:0] out   );//

    always@(*) begin  // This is a combinational circuit
        case(sel)
            0:out = data0;
            1:out = data1;  // begin-end if >1 statement
            2:out = data2;  // begin-end if >1 statement
            3:out = data3;  // begin-end if >1 statement
            4:out =data4;  // begin-end if >1 statement
			5:out = data5;  // begin-end if >1 statement
        default: out = 0;
        endcase
    end

endmodule

//////////////////////////////////////////////////////////////////////////////
//Priority encoder
// synthesis verilog_input_version verilog_2001
module top_module (
    input [3:0] in,
    output reg [1:0] pos  );
	
    always @(*) begin
        case(in)
            4'h0: pos = 2'h0;
			4'h1: pos = 2'h0;
			4'h2: pos = 2'h1;
			4'h3: pos = 2'h0;
			4'h4: pos = 2'h2;
			4'h5: pos = 2'h0;
			4'h6: pos = 2'h1;
			4'h7: pos = 2'h0;
			4'h8: pos = 2'h3;
			4'h9: pos = 2'h0;
			4'ha: pos = 2'h1;
			4'hb: pos = 2'h0;
			4'hc: pos = 2'h2;
			4'hd: pos = 2'h0;
			4'he: pos = 2'h1;
			4'hf: pos = 2'h0;
			default: pos = 2'b0;
        endcase
    end
endmodule

//////////////////////////////////////////////////////////////////////////////
//Priority encoder with casez
// synthesis verilog_input_version verilog_2001
module top_module (
    input [7:0] in,
    output reg [2:0] pos );
    always @(*) begin
        casez (in[7:0])
        8'bzzzzzzz1: pos = 0;   
        8'bzzzzzz1z: pos = 1;
        8'bzzzzz1zz: pos = 2;
        8'bzzzz1zzz: pos = 3;
        8'bzzz1zzzz: pos = 4;   
        8'bzz1zzzzz: pos = 5;
        8'bz1zzzzzz: pos = 6;
        8'b1zzzzzzz: pos = 7;
        
        default: pos = 0;
    	endcase
    end
endmodule
//////////////////////////////////////////////////////////////////////////////
//Avoiding latches
// synthesis verilog_input_version verilog_2001
module top_module (
    input [15:0] scancode,
    output reg left,
    output reg down,
    output reg right,
    output reg up  ); 
    always @(*) begin
        left = 1'b0;	down = 1'b0;  right = 1'b0; 	up = 1'b0;  
        case (scancode)
        16'he06b: left = 1'b1;   
        16'he072: down = ~up; 
        16'he074: right =~left;
        16'he075: up = 1'b1;
    	endcase
    end
endmodule
//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//

//////////////////////////////////////////////////////////////////////////////
//
